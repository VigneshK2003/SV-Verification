-----generator signals-----
 time=0,rst=0,d=1,q=0
-----generator signals-----
 time=0,rst=1,d=0,q=0
-----generator signals-----
 time=0,rst=0,d=0,q=0
-----generator signals-----
 time=0,rst=1,d=0,q=0
-----generator signals-----
 time=0,rst=0,d=1,q=0
--driver signal--
 time=1,rst=0,d=1,q=0
--monitor signals--
 time=5,rst=0,d=1,q=1
--scoreboard signal--
 time=5,rst=0,d=1,q=1
---pass---
--driver signal--
 time=6,rst=1,d=0,q=0
--monitor signals--
 time=10,rst=1,d=0,q=0
--scoreboard signal--
 time=10,rst=1,d=0,q=0
---pass---
--driver signal--
 time=11,rst=0,d=0,q=0
--monitor signals--
 time=15,rst=0,d=0,q=0
--scoreboard signal--
 time=15,rst=0,d=0,q=0
---pass---
--driver signal--
 time=16,rst=1,d=0,q=0
--monitor signals--
 time=20,rst=1,d=0,q=0
--scoreboard signal--
 time=20,rst=1,d=0,q=0
---pass---
--driver signal--
 time=21,rst=0,d=1,q=0
--monitor signals--
 time=25,rst=0,d=1,q=1
--scoreboard signal--
 time=25,rst=0,d=1,q=1
---pass---
$finish at simulation time                   25
           V C S   S i m u l a t i o n   R e p o r t 
