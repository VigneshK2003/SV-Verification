interface intf_df();

   logic clk;
   logic rst;
   logic d;
   logic q;
  
endinterface
