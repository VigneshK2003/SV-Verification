---generator class signals---
time = 0,a = 0,b = 1,c = 1,sum = 0,carry = 0
---generator class signals---
time = 0,a = 1,b = 0,c = 0,sum = 0,carry = 0
---generator class signals---
time = 0,a = 0,b = 0,c = 1,sum = 0,carry = 0
---generator class signals---
time = 0,a = 1,b = 0,c = 0,sum = 0,carry = 0
---generator class signals---
time = 0,a = 0,b = 1,c = 0,sum = 0,carry = 0
---driver signals---
time = 1,a = 0,b = 1,c = 1,sum = 0,carry = 0
---monitor class signal---
time = 5,a = 0,b = 1,c = 1,sum = 0,carry = 1
---signals recieved on scoreboard---
time = 5,a = 0,b = 1,c = 1,sum = 0,carry = 1
------test case passed------
---driver signals---
time = 6,a = 1,b = 0,c = 0,sum = 0,carry = 0
---monitor class signal---
time = 10,a = 1,b = 0,c = 0,sum = 1,carry = 0
---signals recieved on scoreboard---
time = 10,a = 1,b = 0,c = 0,sum = 1,carry = 0
------test case passed------
---driver signals---
time = 11,a = 0,b = 0,c = 1,sum = 0,carry = 0
---monitor class signal---
time = 15,a = 0,b = 0,c = 1,sum = 1,carry = 0
---signals recieved on scoreboard---
time = 15,a = 0,b = 0,c = 1,sum = 1,carry = 0
------test case passed------
---driver signals---
time = 16,a = 1,b = 0,c = 0,sum = 0,carry = 0
---monitor class signal---
time = 20,a = 1,b = 0,c = 0,sum = 1,carry = 0
---signals recieved on scoreboard---
time = 20,a = 1,b = 0,c = 0,sum = 1,carry = 0
------test case passed------
---driver signals---
time = 21,a = 0,b = 1,c = 0,sum = 0,carry = 0
---monitor class signal---
time = 25,a = 0,b = 1,c = 0,sum = 1,carry = 0
---signals recieved on scoreboard---
time = 25,a = 0,b = 1,c = 0,sum = 1,carry = 0
------test case passed------
           V C S   S i m u l a t i o n   R e p o r t 
